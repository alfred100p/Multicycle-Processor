module dec16(ip,clk,i1,i2,i3,i4,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15);
input ip,i1,i2,i3,i4,clk;
output reg o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15;
initial begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end

always@(*)
begin
if(~i1&~i2&~i3&~i4)
begin
o0=ip&clk;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&~i2&~i3&i4)
begin
o0=1'd0;
o1=ip&clk;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&~i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=ip&clk;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&~i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=ip&clk;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&~i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=ip&clk;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&~i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=ip&clk;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=ip&clk;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=ip&clk;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&~i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=ip&clk;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&~i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=ip&clk;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=ip&clk;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=ip&clk;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&i2&~i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=ip&clk;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&i2&~i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=ip&clk;
o14=1'd0;
o15=1'd0;
end
else if(i1&i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=ip&clk;
o15=1'd0;
end
else if(i1&i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=ip&clk;
end
end

endmodule