module dec16(ip,i1,i2,i3,i4,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15);
input ip,i1,i2,i3,i4;
output reg o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15;
initial begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
always@(*)
begin
if(~i1&~i2&~i3&~i4)
begin
o0=1'd1;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&~i2&~i3&i4)
begin
o0=1'd0;
o1=1'd1;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&~i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd1;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&~i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd1;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&~i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd1;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&~i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd1;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd1;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(~i1&i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd1;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&~i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd1;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&~i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd1;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd1;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&~i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd1;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&i2&~i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd1;
o13=1'd0;
o14=1'd0;
o15=1'd0;
end
else if(i1&i2&~i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd1;
o14=1'd0;
o15=1'd0;
end
else if(i1&i2&i3&~i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd1;
o15=1'd0;
end
else if(i1&i2&i3&i4)
begin
o0=1'd0;
o1=1'd0;
o2=1'd0;
o3=1'd0;
o4=1'd0;
o5=1'd0;
o6=1'd0;
o7=1'd0;
o8=1'd0;
o9=1'd0;
o10=1'd0;
o11=1'd0;
o12=1'd0;
o13=1'd0;
o14=1'd0;
o15=1'd1;
end
end

endmodule