`include "dff.v"
module reg16(ip,clk,rst,op);
input [15:0]ip;
input clk,rst;
output [15:0]op;
dff d0(ip[0],clk,rst,op[0]);
dff d1(ip[1],clk,rst,op[1]);
dff d2(ip[2],clk,rst,op[2]);
dff d3(ip[3],clk,rst,op[3]);
dff d4(ip[4],clk,rst,op[4]);
dff d5(ip[5],clk,rst,op[5]);
dff d6(ip[6],clk,rst,op[6]);
dff d7(ip[7],clk,rst,op[7]);
dff d8(ip[8],clk,rst,op[8]);
dff d9(ip[9],clk,rst,op[9]);
dff d10(ip[10],clk,rst,op[10]);
dff d11(ip[11],clk,rst,op[11]);
dff d12(ip[12],clk,rst,op[12]);
dff d13(ip[13],clk,rst,op[13]);
dff d14(ip[14],clk,rst,op[14]);
dff d15(ip[15],clk,rst,op[15]);
endmodule